    `define DATA_WIDTH 16
    `define ADDR_WIDTH 3
    